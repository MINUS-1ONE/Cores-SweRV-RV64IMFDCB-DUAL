// SPDX-License-Identifier: Apache-2.0
// Copyright 2019 Western Digital Corporation or its affiliates.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
package swerv_types;

// used to inst trace, to output dasm info to log file
// performance monitor stuff
typedef struct packed {
                       logic [2:0] trace_rv_i_valid_ip;
                       logic [95:0] trace_rv_i_insn_ip;     //32*3
                       logic [191:0] trace_rv_i_address_ip;  //64*3
                       logic [2:0] trace_rv_i_exception_ip;
                       logic [4:0] trace_rv_i_ecause_ip;    
                       logic [2:0] trace_rv_i_interrupt_ip;
                       logic [63:0] trace_rv_i_tval_ip;     //64
                       } trace_pkt_t;


typedef enum logic [4:0] {
                          NULL      = 5'b00000,
                          MUL       = 5'b00001,
                          LOAD      = 5'b00010,
                          STORE     = 5'b00011,
                          ALU       = 5'b00100,
                          CSRREAD   = 5'b00101,
                          CSRWRITE  = 5'b00110,
                          CSRRW     = 5'b00111,
                          EBREAK    = 5'b01000,
                          ECALL     = 5'b01001,
                          FENCE     = 5'b01010,
                          FENCEI    = 5'b01011,
                          MRET      = 5'b01100,
                          CONDBR    = 5'b01101,
                          JAL       = 5'b01110,
                          BITMANIPU = 5'b01111,
                          ATOMIC    = 5'b10000,
                          LR        = 5'b10001,
                          SC        = 5'b10010
                          } inst_t;

// used to transfer icache data error hamming code info
// because 64bit inst's len is also 32bit, for iacche data bank and error info package we need not any change
typedef struct packed {
`ifdef RV_ICACHE_ECC
                       logic [39:0] ecc;
`else
                       logic [7:0] parity;
`endif
                       } icache_err_pkt_t;

typedef struct packed {
                       logic valid;
                       logic wb;
                       logic [`RV_LSU_NUM_NBLOAD_WIDTH-1:0] tag;
                       logic [4:0] rd;
                       } load_cam_pkt_t;

typedef struct packed {
                       logic pc0_call;
                       logic pc0_ret;
                       logic pc0_pc4;
                       logic pc1_call;
                       logic pc1_ret;
                       logic pc1_pc4;
                       } rets_pkt_t;

// modified prett width from 31 to 63
typedef struct packed {
                       logic valid;
                       logic [11:0] toffset;
                       logic [1:0] hist;
                       logic br_error;
                       logic br_start_error;
                       logic [`RV_BTB_ADDR_HI:`RV_BTB_ADDR_LO] index;
                       logic [1:0] bank;
                       logic [63:1] prett;  // predicted ret target
                       logic [`RV_BHT_GHR_RANGE] fghr;
`ifdef RV_BTB_48
                       logic [1:0] way;
`else
                       logic way;
`endif
                       logic ret;
                       logic [`RV_BTB_BTAG_SIZE-1:0] btag;
                       } br_pkt_t;

typedef struct packed {
                       logic valid;
                       logic [1:0] hist;
                       logic br_error;
                       logic br_start_error;
                       logic [`RV_BTB_ADDR_HI:`RV_BTB_ADDR_LO] index;
                       logic [1:0] bank;
                       logic [`RV_BHT_GHR_RANGE] fghr;
`ifdef RV_BTB_48
                       logic [1:0] way;
`else
                       logic way;
`endif
                       logic middle;
                       } br_tlu_pkt_t;

// modified prett width from 31 to 63
typedef struct packed {
                       logic misp;
                       logic ataken;
                       logic boffset;
                       logic pc4;
                       logic [1:0] hist;
                       logic [11:0] toffset;
                       logic [`RV_BTB_ADDR_HI:`RV_BTB_ADDR_LO] index;
                       logic [1:0] bank;
                       logic valid;
                       logic br_error;
                       logic br_start_error;
                       logic [63:1] prett;
                       logic pcall;
                       logic pret;
                       logic pja;
                       logic [`RV_BTB_BTAG_SIZE-1:0] btag;
                       logic [`RV_BHT_GHR_RANGE] fghr;
`ifdef RV_BTB_48
                       logic [1:0] way;
`else
                       logic way;
`endif
                       } predict_pkt_t;

typedef struct packed {
                       logic legal;
                       logic icaf;
                       logic icaf_second;
                       logic perr;
                       logic sbecc;
                       logic fence_i;
                       logic [3:0] i0trigger;
                       logic [3:0] i1trigger;
                       inst_t pmu_i0_itype;        // pmu - instruction type
                       inst_t pmu_i1_itype;        // pmu - instruction type
                       logic pmu_i0_br_unpred;     // pmu
                       logic pmu_i1_br_unpred;     // pmu
                       logic pmu_divide;
                       logic pmu_lsu_misaligned;
                       } trap_pkt_t;

typedef struct packed {
                       logic [4:0] i0rd;
                       logic i0mul;
                       logic i0load;
                       logic i0store;
                       logic i0div;
                       logic i0v;
                       logic i0valid;
                       logic i0secondary;
                       logic [1:0] i0rs1bype2;
                       logic [1:0] i0rs2bype2;
                       logic [3:0] i0rs1bype3;
                       logic [3:0] i0rs2bype3;
                       logic [4:0] i1rd;
                       logic i1mul;
                       logic i1load;
                       logic i1store;
                       logic i1v;
                       logic i1valid;
                       logic csrwen;
                       logic csrwonly;
                       logic [11:0] csrwaddr;
                       logic i1secondary;
                       logic [1:0] i1rs1bype2;
                       logic [1:0] i1rs2bype2;
                       logic [6:0] i1rs1bype3;
                       logic [6:0] i1rs2bype3;
                       //*******FPU related modify begin******
                       logic i0_fpu;
                       logic i0_wr_frd;
                       logic [4:0] i0_frd;
                       logic i0_fp_to_int;
                       logic i0_int_to_fp;
                       logic i0_fp_to_fp;
                       logic i0_fma;
                       logic fdiv_fsqrt;
                       logic i0_fl;
                       logic i0_fs;
                       logic i1_fpu;
                       logic i1_wr_frd;
                       logic [4:0] i1_frd;
                       logic i1_fp_to_int;
                       logic i1_int_to_fp; 
                       logic i1_fp_to_fp; 
                       logic i1_fma;
                       logic i1_fl;
                       logic i1_fs;
                       //*******FPU related modify end******
                       } dest_pkt_t;

typedef struct packed {
                       logic mul;
                       logic load;
                       logic sec;
                       logic alu;
                       //*******FPU related modify begin******
                       logic fp_to_int;
                       logic int_to_fp;
                       logic fp_to_fp;                       
                       logic fma;
                       logic fl;
                       //*******FPU related modify end******
                       } class_pkt_t;

typedef struct packed {
                       logic [4:0] rs1;
                       logic [4:0] rs2;
                       logic [4:0] rd;
                       //*******FPU related modify begin******
                       logic [4:0] frs1;
                       logic [4:0] frs2;
                       logic [4:0] frs3;
                       logic [4:0] frd;
                       //*******FPU related modify begin******
                       } reg_pkt_t;


typedef struct packed {
                       logic valid;
                       logic land;
                       logic lor;
                       logic lxor;
                       logic sll;
                       logic srl;
                       logic sra;
                       logic beq;
                       logic bne;
                       logic blt;
                       logic bge;
                       logic add;
                       logic sub;
                       logic slt;
                       logic unsign;
                       logic jal;
                       logic predict_t;
                       logic predict_nt;
                       logic csr_write;
                       logic csr_imm;
                       logic word;  // for all alu insts with W-postfix in RV64I

                       // for rvb
                       logic clz;
                       logic ctz;
                       logic cpop;
                       logic sext_b;
                       logic sext_h;
                       logic zext_h;
                       logic min;
                       logic max;
                       logic rol;
                       logic ror;
                       logic bset;
                       logic bclr;
                       logic binv;
                       logic bext;
                       logic sh1add;
                       logic sh2add;
                       logic sh3add;
                       logic orc_b;
                       logic rev8;
                       logic dotuw;
                       logic rs2neg;
                       } alu_pkt_t;

typedef struct packed {
                       logic atomic;
                       logic lr;
                       logic sc;
                       logic [4:0] atomic_instr; // this will be decoded to get which of the amo instruction lsu is doing
                       logic by;
                       logic half;
                       logic word;
                       logic dword;  // for dma and sd/ld inst
                       logic load;
                       logic store;
                       logic unsign;
                       logic dma;    // dma pkt
                       logic store_data_bypass_c1;
                       logic load_ldst_bypass_c1;
                       logic store_data_bypass_c2;
                       logic store_data_bypass_i0_e2_c2;
                       logic [1:0] store_data_bypass_e4_c1;
                       logic [1:0] store_data_bypass_e4_c2;
                       logic [1:0] store_data_bypass_e4_c3;
                       //*******FPU related modify begin******
                       logic fs_data_bypass_c1;
                       logic fs_data_bypass_c2;
                       //*******FPU related modify end******
                       logic valid;
                       } lsu_pkt_t;

typedef struct packed {
                      logic exc_valid;
                      logic single_ecc_error;
                      logic inst_type;   //0: Load, 1: Store
                      logic inst_pipe;   //0: i0, 1: i1
                      logic dma_valid;
                      logic exc_type;    //0: MisAligned, 1: Access Fault
                      logic [63:0] addr;
                      } lsu_error_pkt_t;

typedef struct packed {
                        logic alu;
                        logic rs1;
                        logic rs2;
                        logic imm12;
                        logic rd;
                        logic shimm6;  //adjust from shimm5 to shimm6 for SLLI in RV64I
                        logic imm20;
                        logic pc;
                        logic load;
                        logic store;
                        logic lsu;
                        logic add;
                        logic sub;
                        logic land;
                        logic lor;
                        logic lxor;
                        logic sll;
                        logic sra;
                        logic srl;
                        logic slt;
                        logic unsign;
                        logic condbr;
                        logic beq;
                        logic bne;
                        logic bge;
                        logic blt;
                        logic jal;
                        logic by;
                        logic half;
                        logic word;
                        logic dword;  //added for ld/sd
                        logic csr_read;
                        logic csr_clr;
                        logic csr_set;
                        logic csr_write;
                        logic csr_imm;
                        logic presync;
                        logic postsync;
                        logic ebreak;
                        logic ecall;
                        logic mret;
                        logic mul;
                        logic rs1_sign;
                        logic rs2_sign;
                        logic low;
                        logic div;
                        logic rem;
                        logic fence;
                        logic fence_i;
                        logic pm_alu;
                        logic legal;
                        logic wpostfix;  //for all insts with W-postfix in RV64IM

                        //*******FPU related modify begin******
                        logic fpu;
                        logic frs1; // Need read frs1
                        logic frs2; // Need read frs2
                        logic frs3; // Need read frs3
                        logic frd; // Need write back result to FGPRs
                        logic fflags; // Need write FFLAGS CSR
                        logic fp64;
                        logic islong;
                        logic sign;
                        logic fp_to_int;
                        logic int_to_fp;
                        logic fp_to_fp;
                        logic fma;
                        logic fmin;
                        logic fmax;
                        logic fsgnj;
                        logic fsgnjn;
                        logic fsgnjx;
                        logic fcvt;
                        logic fs;
                        logic fl;
                        logic fclass;
                        logic feq;
                        logic flt;
                        logic fle;
                        logic fmv;
                        logic fadd;
                        logic fsub;
                        logic fmul;
                        logic fmadd;
                        logic fmsub;
                        logic fnmadd;
                        logic fnmsub;
                        logic fdiv;
                        logic fsqrt;
                        //*******FPU related modify end******

                        //for rvb decode
                        logic clz;
                        logic ctz;
                        logic cpop;
                        logic sext_b;
                        logic sext_h;
                        logic zext_h;
                        logic min;
                        logic max;
                        logic rol;
                        logic ror;
                        logic bset;
                        logic bclr;
                        logic binv;
                        logic bext;
                        logic clmul;
                        logic reverse;
                        logic sh1add;
                        logic sh2add;
                        logic sh3add;
                        logic rev8;
                        logic orc_b;
                        logic zba;
                        logic zbb;
                        logic zbc;
                        logic zbs;
                        logic rs2neg;   //for rvb inst that need neg rs2 for example andn/orn/xnor
                        logic dotuw;    //for rvb inst that with .uw postfix for example sh1add.uw/slli.uw
                        logic atomic;
                        logic lr;
                        logic sc;
                       } dec_pkt_t;


typedef struct packed {
                       logic valid;
                       logic rs1_sign;
                       logic rs2_sign;
                       logic word;    //added mulw signal to express MULW inst for RV64M
                       logic low;
                       logic load_mul_rs1_bypass_e1;
                       logic load_mul_rs2_bypass_e1;
                       
                       //added for rvb
                       logic clmul;
                       logic reverse;
                       } mul_pkt_t;

typedef struct packed {
                       logic valid;
                       logic unsign;
                       logic rem;
                       logic word;  //added word signal to express DIV[U]W/REM[U]W inst for RV64M
                       } div_pkt_t;


typedef struct packed {
                        logic        select;
                        logic        match;
                        logic        store;
                        logic        load;
                        logic        execute;
                        logic        m;
                        logic [63:0] tdata2;
            } trigger_pkt_t;


typedef struct packed {
`ifdef RV_ICACHE_ECC
                        logic [74:0]  icache_wrdata; // {dicad1[10:0], dicad0[63:0]}
                                                     // 75 bit for 10 ecc + 32 data
`else
                        logic [65:0]  icache_wrdata; // {dicad0[0:0], dicad0[63:0]}
                                                     // 66 bit for 2 parity + 32 data
`endif
                        logic [18:2]  icache_dicawics;
                        logic         icache_rd_valid;
                        logic         icache_wr_valid;
            } cache_debug_pkt_t;

//******************************************
//*************FPU TYPE START***************
//******************************************
typedef struct packed {
                        logic valid;
                        logic fp_to_int;
                        logic int_to_fp;
                        logic fp_to_fp;
                        logic fma;
                        logic fp64;
                        logic islong;
                        logic sign;
                        logic fmin;
                        logic fmax;
                        logic fsgnj;
                        logic fsgnjn;
                        logic fsgnjx;
                        logic fcvt;
                        logic fs;
                        logic fl;
                        logic fclass;
                        logic feq;
                        logic flt;
                        logic fle;
                        logic fmv;
                        logic fadd;
                        logic fsub;
                        logic fmul;
                        logic fmadd;
                        logic fmsub;
                        logic fnmadd;
                        logic fnmsub;
                        logic fdiv;
                        logic fsqrt;
                        logic [2:0] rm;
                      } fpu_pkt_t;
//******************************************
//*************FPU TYPE END*****************
//******************************************

endpackage // swerv_types
